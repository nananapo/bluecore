package svconfig;
    `ifndef MEMORY_INITIAL_FILE
        `define MEMORY_INITIAL_FILE ""
    `endif
    // メモリの初期値
    localparam MEMORY_INITIAL_FILE = `MEMORY_INITIAL_FILE;
endpackage